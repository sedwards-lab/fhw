`timescale 1ns/1ns
package mMapAdd_package ;
    typedef logic [4:0] \Int4#_t ;
    typedef logic [8:0] \Int8#_t ;
    typedef logic [16:0] \Int16#_t ;
    typedef logic [32:0] \Int#_t ;
    typedef logic [4:0] \Word4#_t ;
    typedef logic [8:0] \Word8#_t ;
    typedef logic [16:0] \Word16#_t ;
    typedef logic [32:0] \Word#_t ;
    typedef logic [5:0] C19_t;
    function C19_t C1_19_dc (logic valid);
      begin
        C1_19_dc = 6'bx;
        C1_19_dc[0:0] = valid;
        C1_19_dc[5:1] = 5'd0;
      end
    endfunction
    function C19_t C2_19_dc (logic valid);
      begin
        C2_19_dc = 6'bx;
        C2_19_dc[0:0] = valid;
        C2_19_dc[5:1] = 5'd1;
      end
    endfunction
    function C19_t C3_19_dc (logic valid);
      begin
        C3_19_dc = 6'bx;
        C3_19_dc[0:0] = valid;
        C3_19_dc[5:1] = 5'd2;
      end
    endfunction
    function C19_t C4_19_dc (logic valid);
      begin
        C4_19_dc = 6'bx;
        C4_19_dc[0:0] = valid;
        C4_19_dc[5:1] = 5'd3;
      end
    endfunction
    function C19_t C5_19_dc (logic valid);
      begin
        C5_19_dc = 6'bx;
        C5_19_dc[0:0] = valid;
        C5_19_dc[5:1] = 5'd4;
      end
    endfunction
    function C19_t C6_19_dc (logic valid);
      begin
        C6_19_dc = 6'bx;
        C6_19_dc[0:0] = valid;
        C6_19_dc[5:1] = 5'd5;
      end
    endfunction
    function C19_t C7_19_dc (logic valid);
      begin
        C7_19_dc = 6'bx;
        C7_19_dc[0:0] = valid;
        C7_19_dc[5:1] = 5'd6;
      end
    endfunction
    function C19_t C8_19_dc (logic valid);
      begin
        C8_19_dc = 6'bx;
        C8_19_dc[0:0] = valid;
        C8_19_dc[5:1] = 5'd7;
      end
    endfunction
    function C19_t C9_19_dc (logic valid);
      begin
        C9_19_dc = 6'bx;
        C9_19_dc[0:0] = valid;
        C9_19_dc[5:1] = 5'd8;
      end
    endfunction
    function C19_t C10_19_dc (logic valid);
      begin
        C10_19_dc = 6'bx;
        C10_19_dc[0:0] = valid;
        C10_19_dc[5:1] = 5'd9;
      end
    endfunction
    function C19_t C11_19_dc (logic valid);
      begin
        C11_19_dc = 6'bx;
        C11_19_dc[0:0] = valid;
        C11_19_dc[5:1] = 5'd10;
      end
    endfunction
    function C19_t C12_19_dc (logic valid);
      begin
        C12_19_dc = 6'bx;
        C12_19_dc[0:0] = valid;
        C12_19_dc[5:1] = 5'd11;
      end
    endfunction
    function C19_t C13_19_dc (logic valid);
      begin
        C13_19_dc = 6'bx;
        C13_19_dc[0:0] = valid;
        C13_19_dc[5:1] = 5'd12;
      end
    endfunction
    function C19_t C14_19_dc (logic valid);
      begin
        C14_19_dc = 6'bx;
        C14_19_dc[0:0] = valid;
        C14_19_dc[5:1] = 5'd13;
      end
    endfunction
    function C19_t C15_19_dc (logic valid);
      begin
        C15_19_dc = 6'bx;
        C15_19_dc[0:0] = valid;
        C15_19_dc[5:1] = 5'd14;
      end
    endfunction
    function C19_t C16_19_dc (logic valid);
      begin
        C16_19_dc = 6'bx;
        C16_19_dc[0:0] = valid;
        C16_19_dc[5:1] = 5'd15;
      end
    endfunction
    function C19_t C17_19_dc (logic valid);
      begin
        C17_19_dc = 6'bx;
        C17_19_dc[0:0] = valid;
        C17_19_dc[5:1] = 5'd16;
      end
    endfunction
    function C19_t C18_19_dc (logic valid);
      begin
        C18_19_dc = 6'bx;
        C18_19_dc[0:0] = valid;
        C18_19_dc[5:1] = 5'd17;
      end
    endfunction
    function C19_t C19_19_dc (logic valid);
      begin
        C19_19_dc = 6'bx;
        C19_19_dc[0:0] = valid;
        C19_19_dc[5:1] = 5'd18;
      end
    endfunction
    typedef logic [1:0] C2_t;
    function C2_t C1_2_dc (logic valid);
      begin
        C1_2_dc = 2'bx;
        C1_2_dc[0:0] = valid;
        C1_2_dc[1:1] = 1'd0;
      end
    endfunction
    function C2_t C2_2_dc (logic valid);
      begin
        C2_2_dc = 2'bx;
        C2_2_dc[0:0] = valid;
        C2_2_dc[1:1] = 1'd1;
      end
    endfunction
    typedef logic [2:0] C3_t;
    function C3_t C1_3_dc (logic valid);
      begin
        C1_3_dc = 3'bx;
        C1_3_dc[0:0] = valid;
        C1_3_dc[2:1] = 2'd0;
      end
    endfunction
    function C3_t C2_3_dc (logic valid);
      begin
        C2_3_dc = 3'bx;
        C2_3_dc[0:0] = valid;
        C2_3_dc[2:1] = 2'd1;
      end
    endfunction
    function C3_t C3_3_dc (logic valid);
      begin
        C3_3_dc = 3'bx;
        C3_3_dc[0:0] = valid;
        C3_3_dc[2:1] = 2'd2;
      end
    endfunction
    typedef logic [0:0] Go_t;
    function Go_t Go_dc (logic valid);
      begin
        Go_dc = 1'bx;
        Go_dc[0:0] = valid;
      end
    endfunction
    typedef logic [16:0] Pointer_QTree_Nat_t;
    function Pointer_QTree_Nat_t Pointer_QTree_Nat_dc (logic valid, \Word16#_t  z1);
      begin
        Pointer_QTree_Nat_dc = 17'bx;
        Pointer_QTree_Nat_dc[0:0] = valid;
        Pointer_QTree_Nat_dc[16:1] = z1[16:1];
      end
    endfunction
    typedef logic [16:0] Pointer_Nat_t;
    function Pointer_Nat_t Pointer_Nat_dc (logic valid, \Word16#_t  z1);
      begin
        Pointer_Nat_dc = 17'bx;
        Pointer_Nat_dc[0:0] = valid;
        Pointer_Nat_dc[16:1] = z1[16:1];
      end
    endfunction
    typedef logic [66:0] QTree_Nat_t;
    function QTree_Nat_t QNone_Nat_dc (logic valid, Go_t z1);
      begin
        QNone_Nat_dc = 67'bx;
        QNone_Nat_dc[0:0] = valid;
        QNone_Nat_dc[2:1] = 2'd0;
        ;
      end
    endfunction
    function QTree_Nat_t QVal_Nat_dc (logic valid, Pointer_Nat_t z1);
      begin
        QVal_Nat_dc = 67'bx;
        QVal_Nat_dc[0:0] = valid;
        QVal_Nat_dc[2:1] = 2'd1;
        QVal_Nat_dc[18:3] = z1[16:1];
      end
    endfunction
    function QTree_Nat_t QNode_Nat_dc (logic valid, Pointer_QTree_Nat_t z1, Pointer_QTree_Nat_t z2, Pointer_QTree_Nat_t z3, Pointer_QTree_Nat_t z4);
      begin
        QNode_Nat_dc = 67'bx;
        QNode_Nat_dc[0:0] = valid;
        QNode_Nat_dc[2:1] = 2'd2;
        QNode_Nat_dc[18:3] = z1[16:1];
        QNode_Nat_dc[34:19] = z2[16:1];
        QNode_Nat_dc[50:35] = z3[16:1];
        QNode_Nat_dc[66:51] = z4[16:1];
      end
    endfunction
    function QTree_Nat_t QError_Nat_dc (logic valid, Go_t z1);
      begin
        QError_Nat_dc = 67'bx;
        QError_Nat_dc[0:0] = valid;
        QError_Nat_dc[2:1] = 2'd3;
        ;
      end
    endfunction
    typedef logic [83:0] MemIn_QTree_Nat_t;
    function MemIn_QTree_Nat_t ReadIn_QTree_Nat_dc (logic valid, \Word16#_t  z1);
      begin
        ReadIn_QTree_Nat_dc = 84'bx;
        ReadIn_QTree_Nat_dc[0:0] = valid;
        ReadIn_QTree_Nat_dc[1:1] = 1'd0;
        ReadIn_QTree_Nat_dc[17:2] = z1[16:1];
      end
    endfunction
    function MemIn_QTree_Nat_t WriteIn_QTree_Nat_dc (logic valid, \Word16#_t  z1, QTree_Nat_t z2);
      begin
        WriteIn_QTree_Nat_dc = 84'bx;
        WriteIn_QTree_Nat_dc[0:0] = valid;
        WriteIn_QTree_Nat_dc[1:1] = 1'd1;
        WriteIn_QTree_Nat_dc[17:2] = z1[16:1];
        WriteIn_QTree_Nat_dc[83:18] = z2[66:1];
      end
    endfunction
    typedef logic [67:0] MemOut_QTree_Nat_t;
    function MemOut_QTree_Nat_t ReadOut_QTree_Nat_dc (logic valid, QTree_Nat_t z1);
      begin
        ReadOut_QTree_Nat_dc = 68'bx;
        ReadOut_QTree_Nat_dc[0:0] = valid;
        ReadOut_QTree_Nat_dc[1:1] = 1'd0;
        ReadOut_QTree_Nat_dc[67:2] = z1[66:1];
      end
    endfunction
    function MemOut_QTree_Nat_t ACK_QTree_Nat_dc (logic valid);
      begin
        ACK_QTree_Nat_dc = 68'bx;
        ACK_QTree_Nat_dc[0:0] = valid;
        ACK_QTree_Nat_dc[1:1] = 1'd1;
      end
    endfunction
    typedef logic [16:0] Pointer_CTf_t;
    function Pointer_CTf_t Pointer_CTf_dc (logic valid, \Word16#_t  z1);
      begin
        Pointer_CTf_dc = 17'bx;
        Pointer_CTf_dc[0:0] = valid;
        Pointer_CTf_dc[16:1] = z1[16:1];
      end
    endfunction
    typedef logic [16:0] Pointer_QTree_Bool_t;
    function Pointer_QTree_Bool_t Pointer_QTree_Bool_dc (logic valid, \Word16#_t  z1);
      begin
        Pointer_QTree_Bool_dc = 17'bx;
        Pointer_QTree_Bool_dc[0:0] = valid;
        Pointer_QTree_Bool_dc[16:1] = z1[16:1];
      end
    endfunction
    typedef logic [115:0] CTf_t;
    function CTf_t Lfsbos_dc (logic valid, Go_t z1);
      begin
        Lfsbos_dc = 116'bx;
        Lfsbos_dc[0:0] = valid;
        Lfsbos_dc[3:1] = 3'd0;
        ;
      end
    endfunction
    function CTf_t Lcall_f3_dc (logic valid, Pointer_CTf_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4, Pointer_QTree_Bool_t z5, Pointer_QTree_Bool_t z6, Pointer_QTree_Bool_t z7);
      begin
        Lcall_f3_dc = 116'bx;
        Lcall_f3_dc[0:0] = valid;
        Lcall_f3_dc[3:1] = 3'd1;
        Lcall_f3_dc[19:4] = z1[16:1];
        Lcall_f3_dc[35:20] = z2[16:1];
        Lcall_f3_dc[51:36] = z3[16:1];
        Lcall_f3_dc[67:52] = z4[16:1];
        Lcall_f3_dc[83:68] = z5[16:1];
        Lcall_f3_dc[99:84] = z6[16:1];
        Lcall_f3_dc[115:100] = z7[16:1];
      end
    endfunction
    function CTf_t Lcall_f2_dc (logic valid, Pointer_QTree_Nat_t z1, Pointer_CTf_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4, Pointer_QTree_Bool_t z5, Pointer_QTree_Bool_t z6);
      begin
        Lcall_f2_dc = 116'bx;
        Lcall_f2_dc[0:0] = valid;
        Lcall_f2_dc[3:1] = 3'd2;
        Lcall_f2_dc[19:4] = z1[16:1];
        Lcall_f2_dc[35:20] = z2[16:1];
        Lcall_f2_dc[51:36] = z3[16:1];
        Lcall_f2_dc[67:52] = z4[16:1];
        Lcall_f2_dc[83:68] = z5[16:1];
        Lcall_f2_dc[99:84] = z6[16:1];
      end
    endfunction
    function CTf_t Lcall_f1_dc (logic valid, Pointer_QTree_Nat_t z1, Pointer_QTree_Nat_t z2, Pointer_CTf_t z3, Pointer_QTree_Bool_t z4, Pointer_QTree_Bool_t z5);
      begin
        Lcall_f1_dc = 116'bx;
        Lcall_f1_dc[0:0] = valid;
        Lcall_f1_dc[3:1] = 3'd3;
        Lcall_f1_dc[19:4] = z1[16:1];
        Lcall_f1_dc[35:20] = z2[16:1];
        Lcall_f1_dc[51:36] = z3[16:1];
        Lcall_f1_dc[67:52] = z4[16:1];
        Lcall_f1_dc[83:68] = z5[16:1];
      end
    endfunction
    function CTf_t Lcall_f0_dc (logic valid, Pointer_QTree_Nat_t z1, Pointer_QTree_Nat_t z2, Pointer_QTree_Nat_t z3, Pointer_CTf_t z4);
      begin
        Lcall_f0_dc = 116'bx;
        Lcall_f0_dc[0:0] = valid;
        Lcall_f0_dc[3:1] = 3'd4;
        Lcall_f0_dc[19:4] = z1[16:1];
        Lcall_f0_dc[35:20] = z2[16:1];
        Lcall_f0_dc[51:36] = z3[16:1];
        Lcall_f0_dc[67:52] = z4[16:1];
      end
    endfunction
    typedef logic [132:0] MemIn_CTf_t;
    function MemIn_CTf_t ReadIn_CTf_dc (logic valid, \Word16#_t  z1);
      begin
        ReadIn_CTf_dc = 133'bx;
        ReadIn_CTf_dc[0:0] = valid;
        ReadIn_CTf_dc[1:1] = 1'd0;
        ReadIn_CTf_dc[17:2] = z1[16:1];
      end
    endfunction
    function MemIn_CTf_t WriteIn_CTf_dc (logic valid, \Word16#_t  z1, CTf_t z2);
      begin
        WriteIn_CTf_dc = 133'bx;
        WriteIn_CTf_dc[0:0] = valid;
        WriteIn_CTf_dc[1:1] = 1'd1;
        WriteIn_CTf_dc[17:2] = z1[16:1];
        WriteIn_CTf_dc[132:18] = z2[115:1];
      end
    endfunction
    typedef logic [116:0] MemOut_CTf_t;
    function MemOut_CTf_t ReadOut_CTf_dc (logic valid, CTf_t z1);
      begin
        ReadOut_CTf_dc = 117'bx;
        ReadOut_CTf_dc[0:0] = valid;
        ReadOut_CTf_dc[1:1] = 1'd0;
        ReadOut_CTf_dc[116:2] = z1[115:1];
      end
    endfunction
    function MemOut_CTf_t ACK_CTf_dc (logic valid);
      begin
        ACK_CTf_dc = 117'bx;
        ACK_CTf_dc[0:0] = valid;
        ACK_CTf_dc[1:1] = 1'd1;
      end
    endfunction
    typedef logic [16:0] \Pointer_CTf''''''''_f''''''''_Bool_t ;
    function \Pointer_CTf''''''''_f''''''''_Bool_t  \Pointer_CTf''''''''_f''''''''_Bool_dc  (logic valid, \Word16#_t  z1);
      begin
        \Pointer_CTf''''''''_f''''''''_Bool_dc  = 17'bx;
        \Pointer_CTf''''''''_f''''''''_Bool_dc [0:0] = valid;
        \Pointer_CTf''''''''_f''''''''_Bool_dc [16:1] = z1[16:1];
      end
    endfunction
    typedef logic [67:0] \CTf''''''''_f''''''''_Bool_t ;
    function \CTf''''''''_f''''''''_Bool_t  \Lf''''''''_f''''''''_Boolsbos_dc  (logic valid, Go_t z1);
      begin
        \Lf''''''''_f''''''''_Boolsbos_dc  = 68'bx;
        \Lf''''''''_f''''''''_Boolsbos_dc [0:0] = valid;
        \Lf''''''''_f''''''''_Boolsbos_dc [3:1] = 3'd0;
        ;
      end
    endfunction
    function \CTf''''''''_f''''''''_Bool_t  \Lcall_f''''''''_f''''''''_Bool3_dc  (logic valid, \Pointer_CTf''''''''_f''''''''_Bool_t  z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4);
      begin
        \Lcall_f''''''''_f''''''''_Bool3_dc  = 68'bx;
        \Lcall_f''''''''_f''''''''_Bool3_dc [0:0] = valid;
        \Lcall_f''''''''_f''''''''_Bool3_dc [3:1] = 3'd1;
        \Lcall_f''''''''_f''''''''_Bool3_dc [19:4] = z1[16:1];
        \Lcall_f''''''''_f''''''''_Bool3_dc [35:20] = z2[16:1];
        \Lcall_f''''''''_f''''''''_Bool3_dc [51:36] = z3[16:1];
        \Lcall_f''''''''_f''''''''_Bool3_dc [67:52] = z4[16:1];
      end
    endfunction
    function \CTf''''''''_f''''''''_Bool_t  \Lcall_f''''''''_f''''''''_Bool2_dc  (logic valid, Pointer_QTree_Nat_t z1, \Pointer_CTf''''''''_f''''''''_Bool_t  z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4);
      begin
        \Lcall_f''''''''_f''''''''_Bool2_dc  = 68'bx;
        \Lcall_f''''''''_f''''''''_Bool2_dc [0:0] = valid;
        \Lcall_f''''''''_f''''''''_Bool2_dc [3:1] = 3'd2;
        \Lcall_f''''''''_f''''''''_Bool2_dc [19:4] = z1[16:1];
        \Lcall_f''''''''_f''''''''_Bool2_dc [35:20] = z2[16:1];
        \Lcall_f''''''''_f''''''''_Bool2_dc [51:36] = z3[16:1];
        \Lcall_f''''''''_f''''''''_Bool2_dc [67:52] = z4[16:1];
      end
    endfunction
    function \CTf''''''''_f''''''''_Bool_t  \Lcall_f''''''''_f''''''''_Bool1_dc  (logic valid, Pointer_QTree_Nat_t z1, Pointer_QTree_Nat_t z2, \Pointer_CTf''''''''_f''''''''_Bool_t  z3, Pointer_QTree_Bool_t z4);
      begin
        \Lcall_f''''''''_f''''''''_Bool1_dc  = 68'bx;
        \Lcall_f''''''''_f''''''''_Bool1_dc [0:0] = valid;
        \Lcall_f''''''''_f''''''''_Bool1_dc [3:1] = 3'd3;
        \Lcall_f''''''''_f''''''''_Bool1_dc [19:4] = z1[16:1];
        \Lcall_f''''''''_f''''''''_Bool1_dc [35:20] = z2[16:1];
        \Lcall_f''''''''_f''''''''_Bool1_dc [51:36] = z3[16:1];
        \Lcall_f''''''''_f''''''''_Bool1_dc [67:52] = z4[16:1];
      end
    endfunction
    function \CTf''''''''_f''''''''_Bool_t  \Lcall_f''''''''_f''''''''_Bool0_dc  (logic valid, Pointer_QTree_Nat_t z1, Pointer_QTree_Nat_t z2, Pointer_QTree_Nat_t z3, \Pointer_CTf''''''''_f''''''''_Bool_t  z4);
      begin
        \Lcall_f''''''''_f''''''''_Bool0_dc  = 68'bx;
        \Lcall_f''''''''_f''''''''_Bool0_dc [0:0] = valid;
        \Lcall_f''''''''_f''''''''_Bool0_dc [3:1] = 3'd4;
        \Lcall_f''''''''_f''''''''_Bool0_dc [19:4] = z1[16:1];
        \Lcall_f''''''''_f''''''''_Bool0_dc [35:20] = z2[16:1];
        \Lcall_f''''''''_f''''''''_Bool0_dc [51:36] = z3[16:1];
        \Lcall_f''''''''_f''''''''_Bool0_dc [67:52] = z4[16:1];
      end
    endfunction
    typedef logic [84:0] \MemIn_CTf''''''''_f''''''''_Bool_t ;
    function \MemIn_CTf''''''''_f''''''''_Bool_t  \ReadIn_CTf''''''''_f''''''''_Bool_dc  (logic valid, \Word16#_t  z1);
      begin
        \ReadIn_CTf''''''''_f''''''''_Bool_dc  = 85'bx;
        \ReadIn_CTf''''''''_f''''''''_Bool_dc [0:0] = valid;
        \ReadIn_CTf''''''''_f''''''''_Bool_dc [1:1] = 1'd0;
        \ReadIn_CTf''''''''_f''''''''_Bool_dc [17:2] = z1[16:1];
      end
    endfunction
    function \MemIn_CTf''''''''_f''''''''_Bool_t  \WriteIn_CTf''''''''_f''''''''_Bool_dc  (logic valid, \Word16#_t  z1, \CTf''''''''_f''''''''_Bool_t  z2);
      begin
        \WriteIn_CTf''''''''_f''''''''_Bool_dc  = 85'bx;
        \WriteIn_CTf''''''''_f''''''''_Bool_dc [0:0] = valid;
        \WriteIn_CTf''''''''_f''''''''_Bool_dc [1:1] = 1'd1;
        \WriteIn_CTf''''''''_f''''''''_Bool_dc [17:2] = z1[16:1];
        \WriteIn_CTf''''''''_f''''''''_Bool_dc [84:18] = z2[67:1];
      end
    endfunction
    typedef logic [68:0] \MemOut_CTf''''''''_f''''''''_Bool_t ;
    function \MemOut_CTf''''''''_f''''''''_Bool_t  \ReadOut_CTf''''''''_f''''''''_Bool_dc  (logic valid, \CTf''''''''_f''''''''_Bool_t  z1);
      begin
        \ReadOut_CTf''''''''_f''''''''_Bool_dc  = 69'bx;
        \ReadOut_CTf''''''''_f''''''''_Bool_dc [0:0] = valid;
        \ReadOut_CTf''''''''_f''''''''_Bool_dc [1:1] = 1'd0;
        \ReadOut_CTf''''''''_f''''''''_Bool_dc [68:2] = z1[67:1];
      end
    endfunction
    function \MemOut_CTf''''''''_f''''''''_Bool_t  \ACK_CTf''''''''_f''''''''_Bool_dc  (logic valid);
      begin
        \ACK_CTf''''''''_f''''''''_Bool_dc  = 69'bx;
        \ACK_CTf''''''''_f''''''''_Bool_dc [0:0] = valid;
        \ACK_CTf''''''''_f''''''''_Bool_dc [1:1] = 1'd1;
      end
    endfunction
    typedef logic [17:0] Nat_t;
    function Nat_t Zero_dc (logic valid, Go_t z1);
      begin
        Zero_dc = 18'bx;
        Zero_dc[0:0] = valid;
        Zero_dc[1:1] = 1'd0;
        ;
      end
    endfunction
    function Nat_t Succ_dc (logic valid, Pointer_Nat_t z1);
      begin
        Succ_dc = 18'bx;
        Succ_dc[0:0] = valid;
        Succ_dc[1:1] = 1'd1;
        Succ_dc[17:2] = z1[16:1];
      end
    endfunction
    typedef logic [34:0] MemIn_Nat_t;
    function MemIn_Nat_t ReadIn_Nat_dc (logic valid, \Word16#_t  z1);
      begin
        ReadIn_Nat_dc = 35'bx;
        ReadIn_Nat_dc[0:0] = valid;
        ReadIn_Nat_dc[1:1] = 1'd0;
        ReadIn_Nat_dc[17:2] = z1[16:1];
      end
    endfunction
    function MemIn_Nat_t WriteIn_Nat_dc (logic valid, \Word16#_t  z1, Nat_t z2);
      begin
        WriteIn_Nat_dc = 35'bx;
        WriteIn_Nat_dc[0:0] = valid;
        WriteIn_Nat_dc[1:1] = 1'd1;
        WriteIn_Nat_dc[17:2] = z1[16:1];
        WriteIn_Nat_dc[34:18] = z2[17:1];
      end
    endfunction
    typedef logic [18:0] MemOut_Nat_t;
    function MemOut_Nat_t ReadOut_Nat_dc (logic valid, Nat_t z1);
      begin
        ReadOut_Nat_dc = 19'bx;
        ReadOut_Nat_dc[0:0] = valid;
        ReadOut_Nat_dc[1:1] = 1'd0;
        ReadOut_Nat_dc[18:2] = z1[17:1];
      end
    endfunction
    function MemOut_Nat_t ACK_Nat_dc (logic valid);
      begin
        ACK_Nat_dc = 19'bx;
        ACK_Nat_dc[0:0] = valid;
        ACK_Nat_dc[1:1] = 1'd1;
      end
    endfunction
    typedef logic [1:0] MyBool_t;
    function MyBool_t MyFalse_dc (logic valid, Go_t z1);
      begin
        MyFalse_dc = 2'bx;
        MyFalse_dc[0:0] = valid;
        MyFalse_dc[1:1] = 1'd0;
        ;
      end
    endfunction
    function MyBool_t MyTrue_dc (logic valid, Go_t z1);
      begin
        MyTrue_dc = 2'bx;
        MyTrue_dc[0:0] = valid;
        MyTrue_dc[1:1] = 1'd1;
        ;
      end
    endfunction
    typedef logic [66:0] QTree_Bool_t;
    function QTree_Bool_t QNone_Bool_dc (logic valid, Go_t z1);
      begin
        QNone_Bool_dc = 67'bx;
        QNone_Bool_dc[0:0] = valid;
        QNone_Bool_dc[2:1] = 2'd0;
        ;
      end
    endfunction
    function QTree_Bool_t QVal_Bool_dc (logic valid, MyBool_t z1);
      begin
        QVal_Bool_dc = 67'bx;
        QVal_Bool_dc[0:0] = valid;
        QVal_Bool_dc[2:1] = 2'd1;
        QVal_Bool_dc[3:3] = z1[1:1];
      end
    endfunction
    function QTree_Bool_t QNode_Bool_dc (logic valid, Pointer_QTree_Bool_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4);
      begin
        QNode_Bool_dc = 67'bx;
        QNode_Bool_dc[0:0] = valid;
        QNode_Bool_dc[2:1] = 2'd2;
        QNode_Bool_dc[18:3] = z1[16:1];
        QNode_Bool_dc[34:19] = z2[16:1];
        QNode_Bool_dc[50:35] = z3[16:1];
        QNode_Bool_dc[66:51] = z4[16:1];
      end
    endfunction
    function QTree_Bool_t QError_Bool_dc (logic valid, Go_t z1);
      begin
        QError_Bool_dc = 67'bx;
        QError_Bool_dc[0:0] = valid;
        QError_Bool_dc[2:1] = 2'd3;
        ;
      end
    endfunction
    typedef logic [83:0] MemIn_QTree_Bool_t;
    function MemIn_QTree_Bool_t ReadIn_QTree_Bool_dc (logic valid, \Word16#_t  z1);
      begin
        ReadIn_QTree_Bool_dc = 84'bx;
        ReadIn_QTree_Bool_dc[0:0] = valid;
        ReadIn_QTree_Bool_dc[1:1] = 1'd0;
        ReadIn_QTree_Bool_dc[17:2] = z1[16:1];
      end
    endfunction
    function MemIn_QTree_Bool_t WriteIn_QTree_Bool_dc (logic valid, \Word16#_t  z1, QTree_Bool_t z2);
      begin
        WriteIn_QTree_Bool_dc = 84'bx;
        WriteIn_QTree_Bool_dc[0:0] = valid;
        WriteIn_QTree_Bool_dc[1:1] = 1'd1;
        WriteIn_QTree_Bool_dc[17:2] = z1[16:1];
        WriteIn_QTree_Bool_dc[83:18] = z2[66:1];
      end
    endfunction
    typedef logic [67:0] MemOut_QTree_Bool_t;
    function MemOut_QTree_Bool_t ReadOut_QTree_Bool_dc (logic valid, QTree_Bool_t z1);
      begin
        ReadOut_QTree_Bool_dc = 68'bx;
        ReadOut_QTree_Bool_dc[0:0] = valid;
        ReadOut_QTree_Bool_dc[1:1] = 1'd0;
        ReadOut_QTree_Bool_dc[67:2] = z1[66:1];
      end
    endfunction
    function MemOut_QTree_Bool_t ACK_QTree_Bool_dc (logic valid);
      begin
        ACK_QTree_Bool_dc = 68'bx;
        ACK_QTree_Bool_dc[0:0] = valid;
        ACK_QTree_Bool_dc[1:1] = 1'd1;
      end
    endfunction
    typedef logic [3:0] C8_t;
    function C8_t C1_8_dc (logic valid);
      begin
        C1_8_dc = 4'bx;
        C1_8_dc[0:0] = valid;
        C1_8_dc[3:1] = 3'd0;
      end
    endfunction
    function C8_t C2_8_dc (logic valid);
      begin
        C2_8_dc = 4'bx;
        C2_8_dc[0:0] = valid;
        C2_8_dc[3:1] = 3'd1;
      end
    endfunction
    function C8_t C3_8_dc (logic valid);
      begin
        C3_8_dc = 4'bx;
        C3_8_dc[0:0] = valid;
        C3_8_dc[3:1] = 3'd2;
      end
    endfunction
    function C8_t C4_8_dc (logic valid);
      begin
        C4_8_dc = 4'bx;
        C4_8_dc[0:0] = valid;
        C4_8_dc[3:1] = 3'd3;
      end
    endfunction
    function C8_t C5_8_dc (logic valid);
      begin
        C5_8_dc = 4'bx;
        C5_8_dc[0:0] = valid;
        C5_8_dc[3:1] = 3'd4;
      end
    endfunction
    function C8_t C6_8_dc (logic valid);
      begin
        C6_8_dc = 4'bx;
        C6_8_dc[0:0] = valid;
        C6_8_dc[3:1] = 3'd5;
      end
    endfunction
    function C8_t C7_8_dc (logic valid);
      begin
        C7_8_dc = 4'bx;
        C7_8_dc[0:0] = valid;
        C7_8_dc[3:1] = 3'd6;
      end
    endfunction
    function C8_t C8_8_dc (logic valid);
      begin
        C8_8_dc = 4'bx;
        C8_8_dc[0:0] = valid;
        C8_8_dc[3:1] = 3'd7;
      end
    endfunction
    typedef logic [4:0] C15_t;
    function C15_t C1_15_dc (logic valid);
      begin
        C1_15_dc = 5'bx;
        C1_15_dc[0:0] = valid;
        C1_15_dc[4:1] = 4'd0;
      end
    endfunction
    function C15_t C2_15_dc (logic valid);
      begin
        C2_15_dc = 5'bx;
        C2_15_dc[0:0] = valid;
        C2_15_dc[4:1] = 4'd1;
      end
    endfunction
    function C15_t C3_15_dc (logic valid);
      begin
        C3_15_dc = 5'bx;
        C3_15_dc[0:0] = valid;
        C3_15_dc[4:1] = 4'd2;
      end
    endfunction
    function C15_t C4_15_dc (logic valid);
      begin
        C4_15_dc = 5'bx;
        C4_15_dc[0:0] = valid;
        C4_15_dc[4:1] = 4'd3;
      end
    endfunction
    function C15_t C5_15_dc (logic valid);
      begin
        C5_15_dc = 5'bx;
        C5_15_dc[0:0] = valid;
        C5_15_dc[4:1] = 4'd4;
      end
    endfunction
    function C15_t C6_15_dc (logic valid);
      begin
        C6_15_dc = 5'bx;
        C6_15_dc[0:0] = valid;
        C6_15_dc[4:1] = 4'd5;
      end
    endfunction
    function C15_t C7_15_dc (logic valid);
      begin
        C7_15_dc = 5'bx;
        C7_15_dc[0:0] = valid;
        C7_15_dc[4:1] = 4'd6;
      end
    endfunction
    function C15_t C8_15_dc (logic valid);
      begin
        C8_15_dc = 5'bx;
        C8_15_dc[0:0] = valid;
        C8_15_dc[4:1] = 4'd7;
      end
    endfunction
    function C15_t C9_15_dc (logic valid);
      begin
        C9_15_dc = 5'bx;
        C9_15_dc[0:0] = valid;
        C9_15_dc[4:1] = 4'd8;
      end
    endfunction
    function C15_t C10_15_dc (logic valid);
      begin
        C10_15_dc = 5'bx;
        C10_15_dc[0:0] = valid;
        C10_15_dc[4:1] = 4'd9;
      end
    endfunction
    function C15_t C11_15_dc (logic valid);
      begin
        C11_15_dc = 5'bx;
        C11_15_dc[0:0] = valid;
        C11_15_dc[4:1] = 4'd10;
      end
    endfunction
    function C15_t C12_15_dc (logic valid);
      begin
        C12_15_dc = 5'bx;
        C12_15_dc[0:0] = valid;
        C12_15_dc[4:1] = 4'd11;
      end
    endfunction
    function C15_t C13_15_dc (logic valid);
      begin
        C13_15_dc = 5'bx;
        C13_15_dc[0:0] = valid;
        C13_15_dc[4:1] = 4'd12;
      end
    endfunction
    function C15_t C14_15_dc (logic valid);
      begin
        C14_15_dc = 5'bx;
        C14_15_dc[0:0] = valid;
        C14_15_dc[4:1] = 4'd13;
      end
    endfunction
    function C15_t C15_15_dc (logic valid);
      begin
        C15_15_dc = 5'bx;
        C15_15_dc[0:0] = valid;
        C15_15_dc[4:1] = 4'd14;
      end
    endfunction
    typedef logic [2:0] C4_t;
    function C4_t C1_4_dc (logic valid);
      begin
        C1_4_dc = 3'bx;
        C1_4_dc[0:0] = valid;
        C1_4_dc[2:1] = 2'd0;
      end
    endfunction
    function C4_t C2_4_dc (logic valid);
      begin
        C2_4_dc = 3'bx;
        C2_4_dc[0:0] = valid;
        C2_4_dc[2:1] = 2'd1;
      end
    endfunction
    function C4_t C3_4_dc (logic valid);
      begin
        C3_4_dc = 3'bx;
        C3_4_dc[0:0] = valid;
        C3_4_dc[2:1] = 2'd2;
      end
    endfunction
    function C4_t C4_4_dc (logic valid);
      begin
        C4_4_dc = 3'bx;
        C4_4_dc[0:0] = valid;
        C4_4_dc[2:1] = 2'd3;
      end
    endfunction
    typedef logic [3:0] C5_t;
    function C5_t C1_5_dc (logic valid);
      begin
        C1_5_dc = 4'bx;
        C1_5_dc[0:0] = valid;
        C1_5_dc[3:1] = 3'd0;
      end
    endfunction
    function C5_t C2_5_dc (logic valid);
      begin
        C2_5_dc = 4'bx;
        C2_5_dc[0:0] = valid;
        C2_5_dc[3:1] = 3'd1;
      end
    endfunction
    function C5_t C3_5_dc (logic valid);
      begin
        C3_5_dc = 4'bx;
        C3_5_dc[0:0] = valid;
        C3_5_dc[3:1] = 3'd2;
      end
    endfunction
    function C5_t C4_5_dc (logic valid);
      begin
        C4_5_dc = 4'bx;
        C4_5_dc[0:0] = valid;
        C4_5_dc[3:1] = 3'd3;
      end
    endfunction
    function C5_t C5_5_dc (logic valid);
      begin
        C5_5_dc = 4'bx;
        C5_5_dc[0:0] = valid;
        C5_5_dc[3:1] = 3'd4;
      end
    endfunction
    typedef logic [32:0] \TupGo___Pointer_QTree_Bool___Pointer_CTf''''''''_f''''''''_Bool_t ;
    function \TupGo___Pointer_QTree_Bool___Pointer_CTf''''''''_f''''''''_Bool_t  \TupGo___Pointer_QTree_Bool___Pointer_CTf''''''''_f''''''''_Bool_dc  (logic valid, Go_t z1, Pointer_QTree_Bool_t z2, \Pointer_CTf''''''''_f''''''''_Bool_t  z3);
      begin
        \TupGo___Pointer_QTree_Bool___Pointer_CTf''''''''_f''''''''_Bool_dc  = 33'bx;
        \TupGo___Pointer_QTree_Bool___Pointer_CTf''''''''_f''''''''_Bool_dc [0:0] = valid;
        ;
        \TupGo___Pointer_QTree_Bool___Pointer_CTf''''''''_f''''''''_Bool_dc [16:1] = z2[16:1];
        \TupGo___Pointer_QTree_Bool___Pointer_CTf''''''''_f''''''''_Bool_dc [32:17] = z3[16:1];
      end
    endfunction
    typedef logic [48:0] TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_t;
    function TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_t TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc (logic valid, Go_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, Pointer_CTf_t z4);
      begin
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc = 49'bx;
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc[0:0] = valid;
        ;
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc[16:1] = z2[16:1];
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc[32:17] = z3[16:1];
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc[48:33] = z4[16:1];
      end
    endfunction
    typedef logic [16:0] TupGo___Pointer_QTree_Bool_t;
    function TupGo___Pointer_QTree_Bool_t TupGo___Pointer_QTree_Bool_dc (logic valid, Go_t z1, Pointer_QTree_Bool_t z2);
      begin
        TupGo___Pointer_QTree_Bool_dc = 17'bx;
        TupGo___Pointer_QTree_Bool_dc[0:0] = valid;
        ;
        TupGo___Pointer_QTree_Bool_dc[16:1] = z2[16:1];
      end
    endfunction
    typedef logic [32:0] TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t;
    function TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc (logic valid, Go_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3);
      begin
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc = 33'bx;
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[0:0] = valid;
        ;
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[16:1] = z2[16:1];
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[32:17] = z3[16:1];
      end
    endfunction
    typedef logic [0:0] TupGo_t;
    function TupGo_t TupGo_dc (logic valid, Go_t z1);
      begin
        TupGo_dc = 1'bx;
        TupGo_dc[0:0] = valid;
        ;
      end
    endfunction
endpackage